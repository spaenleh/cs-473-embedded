
module system (
	clk_clk,
	pwm_out_conduit,
	reset_reset_n);	

	input		clk_clk;
	output		pwm_out_conduit;
	input		reset_reset_n;
endmodule
