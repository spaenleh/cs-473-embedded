
module system (
	clk_clk,
	reset_reset_n,
	parallel_port_export);	

	input		clk_clk;
	input		reset_reset_n;
	inout	[7:0]	parallel_port_export;
endmodule
